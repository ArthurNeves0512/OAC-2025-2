`ifndef PARAM
    `include "Parametros.v"
`endif

module reg_ID_EX (
    input wire clk,
    input wire reset,
    input wire flush,
    
    // id
    input wire [31:0] pc_plus_4_in,
    input wire [31:0] read_data1_in,
    input wire [31:0] read_data2_in,
    input wire [31:0] imm_in,
    input wire [4:0] rs1_in,
    input wire [4:0] rs2_in,
    input wire [4:0] rd_in,
    
    // controle
    input wire ALUSrc_in,
    input wire [1:0] ALUOp_in,
    input wire MemRead_in,
    input wire MemWrite_in,
    input wire Branch_in,
    input wire RegWrite_in,
    input wire MemToReg_in,
    
    // ex
    output reg [31:0] pc_plus_4_out,
    output reg [31:0] read_data1_out,
    output reg [31:0] read_data2_out,
    output reg [31:0] imm_out,
    output reg [4:0] rs1_out,
    output reg [4:0] rs2_out,
    output reg [4:0] rd_out,
    
    output reg ALUSrc_out,
    output reg [1:0] ALUOp_out,
    output reg MemRead_out,
    output reg MemWrite_out,
    output reg Branch_out,
    output reg RegWrite_out,
    output reg MemToReg_out
);

    always @(posedge clk or posedge reset) begin
        if (reset || flush) begin
            pc_plus_4_out <= 32'b0;
            read_data1_out <= 32'b0;
            read_data2_out <= 32'b0;
            imm_out <= 32'b0;
            rs1_out <= 5'b0;
            rs2_out <= 5'b0;
            rd_out <= 5'b0;
            ALUSrc_out <= 1'b0;
            ALUOp_out <= 2'b0;
            MemRead_out <= 1'b0;
            MemWrite_out <= 1'b0;
            Branch_out <= 1'b0;
            RegWrite_out <= 1'b0;
            MemToReg_out <= 1'b0;
        end else begin
            pc_plus_4_out <= pc_plus_4_in;
            read_data1_out <= read_data1_in;
            read_data2_out <= read_data2_in;
            imm_out <= imm_in;
            rs1_out <= rs1_in;
            rs2_out <= rs2_in;
            rd_out <= rd_in;
            ALUSrc_out <= ALUSrc_in;
            ALUOp_out <= ALUOp_in;
            MemRead_out <= MemRead_in;
            MemWrite_out <= MemWrite_in;
            Branch_out <= Branch_in;
            RegWrite_out <= RegWrite_in;
            MemToReg_out <= MemToReg_in;
        end
    end

endmodule